`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2021  Matthew J. Dovey
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <https://www.gnu.org/licenses/>.
// 
// Create Date: 01.12.2021 20:40:15
// Module Name: resets
// 
//////////////////////////////////////////////////////////////////////////////////


module audio_reset (
(* X_INTERFACE_PARAMETER = "POLARITY ACTIVE_LOW" *)  
    input   resetn,
    
(* X_INTERFACE_PARAMETER = "POLARITY ACTIVE_HIGH" *)  
(* ASYNC_REG = "TRUE" *)
    output reg rst,

(* X_INTERFACE_PARAMETER = "POLARITY ACTIVE_LOW" *)  
(* ASYNC_REG = "TRUE" *)
    output reg rstn,

(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 clk CLK" *)
(* X_INTERFACE_PARAMETER = "ASSOCIATED_RESET rst:rstn" *)
    input clk
);
    
    always @(posedge clk)
    begin
        rst  <= ~resetn;
        rstn <=  resetn;
    end
    
endmodule

